.subckt ideal_diode a k Vf=0.7
* Subcircuit Body
	s1 a ki a ki mysw
	c1 a k 0.1n
	vdiode ki k {Vf}
	.model mysw sw vt=0 vh=0 ron=1e-3 roff=1e7
.ends name